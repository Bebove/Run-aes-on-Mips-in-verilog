`timescale 1 ns / 1 ps 
module Instruction_memory (reset,addr,rd);
  input reset;
  input[31:0]  addr;
  output[31:0]  rd;
  reg[31:0]   RAM[255:0];
  assign rd = RAM[addr[31:2]];
  
  always@(negedge reset)
  begin
//keygen part
RAM[ 0]<=32'b001000_00000_00001_00000_100010110_00; //addi 278->reg1
RAM[ 1]<=32'b001000_00000_11101_00000_111000100_00; //addi 452*4->reg29
RAM[ 2]<=32'b001000_00000_11100_00000_111001110_00; //addi 462*4->reg28
RAM[ 3]<=32'b001000_00000_11111_00000_100010011_01; //addi 275->reg31

//FIRST_ROW
RAM[ 4]<=32'b100011_00001_00010_00000_000000100_00; //lw +4 reg2
RAM[ 5]<=32'b100011_00001_00011_00000_000001000_00; //lw +8 reg3
RAM[ 6]<=32'b100011_00001_00100_00000_000001100_00; //lw +12 reg4 
RAM[ 7]<=32'b100011_00001_00101_00000_000000000_00; //lw +0 reg5
RAM[ 8]<=32'b000000_00000_00010_00010_00010_000000; //reg2 <<2
RAM[ 9]<=32'b000000_00000_00011_00011_00010_000000; //reg3 <<2
RAM[10]<=32'b000000_00000_00100_00100_00010_000000; //reg4 <<2
RAM[11]<=32'b000000_00000_00101_00101_00010_000000; //reg5 <<2
RAM[12]<=32'b100011_00010_00110_00000_000000000_00; //lw  reg2 reg6
RAM[13]<=32'b100011_00011_00111_00000_000000000_00; //lw  reg3 reg7
RAM[14]<=32'b100011_00100_01000_00000_000000000_00; //lw  reg4 reg8
RAM[15]<=32'b100011_00101_01001_00000_000000000_00; //lw  reg5 reg9
RAM[16]<=32'b100011_11101_11110_00000_000000000_00; //lw reg29 reg30
RAM[17]<=32'b001000_11101_11101_00000_000000001_00; //addi  reg29 + 4
RAM[18]<=32'b000000_00110_11110_00110_00000_100110; //xor
RAM[19]<=32'b000000_00111_00000_00111_00000_100110; //xor
RAM[20]<=32'b000000_01000_00000_01000_00000_100110; //xor
RAM[21]<=32'b000000_01001_00000_01001_00000_100110; //xor
RAM[22]<=32'b100011_11111_00101_00000_000000000_00; //lw +0 reg2
RAM[23]<=32'b100011_11111_00010_00000_000000100_00; //lw +4 reg3
RAM[24]<=32'b100011_11111_00011_00000_000001000_00; //lw +8 reg4
RAM[25]<=32'b100011_11111_00100_00000_000001100_00; //lw +12 reg5 
RAM[26]<=32'b000000_00110_00101_00110_00000_100110; //xor
RAM[27]<=32'b000000_00111_00010_00111_00000_100110; //xor
RAM[28]<=32'b000000_01000_00011_01000_00000_100110; //xor
RAM[29]<=32'b000000_01001_00100_01001_00000_100110; //xor
RAM[30]<=32'b101011_00001_00110_00000_000001101_00; //sw +13
RAM[31]<=32'b101011_00001_00111_00000_000010001_00; //sw +13+4
RAM[32]<=32'b101011_00001_01000_00000_000010101_00; //sw +13+8
RAM[33]<=32'b101011_00001_01001_00000_000011001_00; //sw +13+12

RAM[34]<=32'b001000_11111_11111_00000_000000001_00; //addi reg31+4->reg31
RAM[35]<=32'b100011_11111_00101_00000_000000000_00; //lw +0 reg2
RAM[36]<=32'b100011_11111_00010_00000_000000100_00; //lw +4 reg3
RAM[37]<=32'b100011_11111_00011_00000_000001000_00; //lw +8 reg4
RAM[38]<=32'b100011_11111_00100_00000_000001100_00; //lw +12 reg5 
RAM[39]<=32'b000000_00110_00101_00110_00000_100110; //xor
RAM[40]<=32'b000000_00111_00010_00111_00000_100110; //xor
RAM[41]<=32'b000000_01000_00011_01000_00000_100110; //xor
RAM[42]<=32'b000000_01001_00100_01001_00000_100110; //xor
RAM[43]<=32'b101011_00001_00110_00000_000001110_00; //sw +13+1
RAM[44]<=32'b101011_00001_00111_00000_000010010_00; //sw +13+4+1
RAM[45]<=32'b101011_00001_01000_00000_000010110_00; //sw +13+8+1
RAM[46]<=32'b101011_00001_01001_00000_000011010_00; //sw +13+12+1

RAM[47]<=32'b001000_11111_11111_00000_000000001_00; //addi reg31+4->reg31
RAM[48]<=32'b100011_11111_00101_00000_000000000_00; //lw +0 reg2
RAM[49]<=32'b100011_11111_00010_00000_000000100_00; //lw +4 reg3
RAM[50]<=32'b100011_11111_00011_00000_000001000_00; //lw +8 reg4
RAM[51]<=32'b100011_11111_00100_00000_000001100_00; //lw +12 reg5 
RAM[52]<=32'b000000_00110_00101_00110_00000_100110; //xor
RAM[53]<=32'b000000_00111_00010_00111_00000_100110; //xor
RAM[54]<=32'b000000_01000_00011_01000_00000_100110; //xor
RAM[55]<=32'b000000_01001_00100_01001_00000_100110; //xor
RAM[56]<=32'b101011_00001_00110_00000_000001111_00; //sw +13+2
RAM[57]<=32'b101011_00001_00111_00000_000010011_00; //sw +13+4+2
RAM[58]<=32'b101011_00001_01000_00000_000010111_00; //sw +13+8+2
RAM[59]<=32'b101011_00001_01001_00000_000011011_00; //sw +13+12+2


RAM[60]<=32'b001000_11111_11111_00000_000000001_00; //addi reg31+4->reg31
RAM[61]<=32'b100011_11111_00101_00000_000000000_00; //lw +0 reg2
RAM[62]<=32'b100011_11111_00010_00000_000000100_00; //lw +4 reg3
RAM[63]<=32'b100011_11111_00011_00000_000001000_00; //lw +8 reg4
RAM[64]<=32'b100011_11111_00100_00000_000001100_00; //lw +12 reg5 
RAM[65]<=32'b000000_00110_00101_00110_00000_100110; //xor
RAM[66]<=32'b000000_00111_00010_00111_00000_100110; //xor
RAM[67]<=32'b000000_01000_00011_01000_00000_100110; //xor
RAM[68]<=32'b000000_01001_00100_01001_00000_100110; //xor
RAM[69]<=32'b101011_00001_00110_00000_000010000_00; //sw +13+3
RAM[70]<=32'b101011_00001_00111_00000_000010100_00; //sw +13+4+3
RAM[71]<=32'b101011_00001_01000_00000_000011000_00; //sw +13+8+3
RAM[72]<=32'b101011_00001_01001_00000_000011100_00; //sw +13+12+3
//FIRST_ROW done
RAM[73]<=32'b001000_11111_11111_00000_000001101_00; //addi reg31+13->reg31
RAM[74]<=32'b001000_00001_00001_00000_000010000_00; //update reg1 + 16
RAM[75]<=32'b000101_11101_11100_11111_110111000_00; //bne reg29==��ֹ��ַreg28? continue:pc-72*4







//aes part
//Addroundkey(use reg20 reg21 reg22 reg 16 reg17,fuse reg25)
RAM[76]<=32'b100011_00000_10100_00000_111000011_00; //lw data[451).initial=275->reg20
RAM[77]<=32'b100011_00000_10101_00000_100000010_00; //lw data[258)=259->reg21
RAM[78]<=32'b001000_10101_11001_00000_000010000_00; //addi 259+16 =275->reg25
RAM[79]<=32'b001000_10101_11110_00000_000000001_00; //addi copy to 11110
RAM[80]<=32'b100011_10100_10110_00000_000000000_00; //lw 
RAM[81]<=32'b100011_10101_10000_00000_000000000_00; //lw
RAM[82]<=32'b000000_10110_10000_10001_00000_100110; //xor
RAM[83]<=32'b101011_10101_10001_00000_000000000_00; //sw
RAM[84]<=32'b001000_10100_10100_00000_000000001_00; //addi
RAM[85]<=32'b001000_10101_10101_00000_000000001_00; //addi
RAM[86]<=32'b000101_11110_11001_11111_111111000_00; //bne reg21==reg25? continue:pc-7*4
RAM[87]<=32'b101011_00000_10100_00000_111000011_00; //sw reg20->data[451)


//the BIGround begin ,use reg23 24 as counter
RAM[88]<=32'b001000_00000_11000_00000_000000010_10; //addi set counter n to reg 24
RAM[89]<=32'b001000_00000_10111_00000_000000000_00; //addi set 0 to reg 23
//BIGround bnepoint
RAM[90]<=32'b001000_10111_10111_00000_000000000_01; //set 23=23+1
//subbyte(use reg21 reg2 reg3, fuse reg25)
RAM[91]<=32'b100011_00000_10101_00000_100000010_00; //lw lw data[258)=259->reg21
RAM[92]<=32'b100011_10101_00010_00000_000000000_00; //lw data to reg2
RAM[93]<=32'b000000_00000_00010_00010_00010_000000; //reg2 <<2
RAM[94]<=32'b001000_10101_11110_00000_000000001_00; //addi reg21 copy to 11110
RAM[95]<=32'b100011_00010_00011_00000_000000000_00; //lw the sbox code to reg3
RAM[96]<=32'b101011_10101_00011_00000_000000000_00; //sw reg3 to data
RAM[97]<=32'b001000_10101_10101_00000_000000001_00; //addi reg21
RAM[98]<=32'b000101_11110_11001_11111_111111001_00; //bne reg21==reg25? continue:pc-7*4

//ShiftRows(use reg5-16)
RAM[99]<=32'b100011_00000_00101_00000_100000111_00; //lw data to reg5
RAM[100]<=32'b100011_00000_00110_00000_100001000_00; //lw data to reg6
RAM[101]<=32'b100011_00000_00111_00000_100001001_00; //lw data to reg7
RAM[102]<=32'b100011_00000_01000_00000_100001010_00; //lw data to reg8
RAM[103]<=32'b100011_00000_01001_00000_100001011_00; //lw data to reg9
RAM[104]<=32'b100011_00000_01010_00000_100001100_00; //lw data to reg10
RAM[105]<=32'b100011_00000_01011_00000_100001101_00; //lw data to reg11
RAM[106]<=32'b100011_00000_01100_00000_100001110_00; //lw data to reg12
RAM[107]<=32'b100011_00000_01101_00000_100001111_00; //lw data to reg13
RAM[108]<=32'b100011_00000_01110_00000_100010000_00; //lw data to reg14
RAM[109]<=32'b100011_00000_01111_00000_100010001_00; //lw data to reg15
RAM[110]<=32'b100011_00000_10000_00000_100010010_00; //lw data to reg16
RAM[111]<=32'b101011_00000_00110_00000_100000111_00; //sw data from reg6
RAM[112]<=32'b101011_00000_00111_00000_100001000_00; //sw data from reg7
RAM[113]<=32'b101011_00000_01000_00000_100001001_00; //sw data from reg8
RAM[114]<=32'b101011_00000_00101_00000_100001010_00; //sw data from reg5
RAM[115]<=32'b101011_00000_01011_00000_100001011_00; //sw data from reg11
RAM[116]<=32'b101011_00000_01100_00000_100001100_00; //sw data from reg12
RAM[117]<=32'b101011_00000_01001_00000_100001101_00; //sw data from reg9
RAM[118]<=32'b101011_00000_01010_00000_100001110_00; //sw data from reg10
RAM[119]<=32'b101011_00000_10000_00000_100001111_00; //sw data from reg16
RAM[120]<=32'b101011_00000_01101_00000_100010000_00; //sw data from reg13
RAM[121]<=32'b101011_00000_01110_00000_100010001_00; //sw data from reg14
RAM[122]<=32'b101011_00000_01111_00000_100010010_00; //sw data from reg15
//the bne for the last round of BIGround
RAM[123]<=32'b000100_11000_10111_00000_000110101_00; //beq reg23==reg24? pc-99*4:continue
//Mixcolumns:
//  fixreg:30 29 28 27 26 31;
//  data_reg:2,3,4,5;
//  2_reg :7,8,9,10;
//  3_reg :11,12,13,14;
//  xor_reg :15,16,17,18;
//compare_reg:19,20,21,22; 
RAM[124]<=32'b001000_00000_11110_00000_0000111_1111; //addi reg0 0111_1111 reg30 �Ƚϳ���
RAM[125]<=32'b001000_00000_11101_00000_0000000_0001; //addi reg0 0000_0001 reg29 1����
RAM[126]<=32'b001000_00000_11100_00000_0000001_1011; //addi reg0 0001_1011 reg28 xor����
RAM[127]<=32'b100011_00000_11011_00000_100000010_00; //lw  data[258)=259-> reg27 ���ݳ�ʼ��ַ
RAM[128]<=32'b100011_00000_11010_00000_100000010_00; //lw   ����һ�ݵ�ַ��reg26
RAM[129]<=32'b001000_11010_11111_00000_000000100_00; //addi ������ֹ��ַreg26+4��reg31
//load �����ݵ�reg2��3��4��5,����λ����
RAM[130]<=32'b100011_11011_00010_00000_000000000_00; //lw data[reg21+0)   reg2
RAM[131]<=32'b100011_11011_00011_00000_000000100_00; //lw data[reg21+4)   reg3
RAM[132]<=32'b100011_11011_00100_00000_000001000_00; //lw data[reg21+8)   reg4
RAM[133]<=32'b100011_11011_00101_00000_000001100_00; //lw data[reg21+12)  reg5
RAM[134]<=32'b000000_00000_00010_00111_11001_000000; //ͳһ��λreg2->reg7
RAM[135]<=32'b000000_00000_00011_01000_11001_000000; //ͳһ��λreg3->reg8
RAM[136]<=32'b000000_00000_00100_01001_11001_000000; //ͳһ��λreg4->reg9
RAM[137]<=32'b000000_00000_00101_01010_11001_000000; //ͳһ��λreg5->reg10
RAM[138]<=32'b000000_00000_00111_00111_11000_000010; //ͳһ��λreg7->reg7
RAM[139]<=32'b000000_00000_01000_01000_11000_000010; //ͳһ��λreg8->reg8
RAM[140]<=32'b000000_00000_01001_01001_11000_000010; //ͳһ��λreg9->reg9
RAM[141]<=32'b000000_00000_01010_01010_11000_000010; //ͳһ��λreg10->reg10
//data_compare
RAM[142]<=32'b000000_11110_00010_10011_00000_101010; //slt reg30reg2reg19 �ж������Ƿ��?0111_1111��,����ڰ�λ�?1������Ҫ���?
RAM[143]<=32'b000000_11110_00011_10100_00000_101010; //slt reg30reg3reg20 �ж������Ƿ��?0111_1111��,����ڰ�λ�?1������Ҫ���?
RAM[144]<=32'b000000_11110_00100_10101_00000_101010; //slt reg30reg4reg21 �ж������Ƿ��?0111_1111��,����ڰ�λ�?1������Ҫ���?
RAM[145]<=32'b000000_11110_00101_10110_00000_101010; //slt reg30reg5reg22 �ж������Ƿ��?0111_1111��,����ڰ�λ�?1������Ҫ���?
//data1
RAM[146]<=32'b000101_10011_11101_00000_000000001_00; //bne reg6 1  pc+4+4  //reg6=0!=1,����Ҫ����������ת
RAM[147]<=32'b000000_11100_00111_00111_00000_100110; //����ת����==1����˵��Ҫ����xor��reg7��
RAM[148]<=32'b000000_00010_00111_01011_00000_100110; //������ת��񣬶�Ҫ��s����xor��reg11��
//data2
RAM[149]<=32'b000101_10100_11101_00000_000000001_00; 
RAM[150]<=32'b000000_11100_01000_01000_00000_100110; //reg8 
RAM[151]<=32'b000000_00011_01000_01100_00000_100110; //reg12
//data3
RAM[152]<=32'b000101_10101_11101_00000_000000001_00; 
RAM[153]<=32'b000000_11100_01001_01001_00000_100110; //reg9
RAM[154]<=32'b000000_00100_01001_01101_00000_100110; //reg13
//data4
RAM[155]<=32'b000101_10110_11101_00000_000000001_00; 
RAM[156]<=32'b000000_11100_01010_01010_00000_100110; //reg10
RAM[157]<=32'b000000_00101_01010_01110_00000_100110; //reg14
//xor reg7 reg12 reg4 reg5 =>reg15
RAM[158]<=32'b000000_00111_01100_01111_00000_100110;
RAM[159]<=32'b000000_00100_01111_01111_00000_100110;
RAM[160]<=32'b000000_00101_01111_01111_00000_100110;
//xor reg2 reg8  reg13 reg5 =>reg16
RAM[161]<=32'b000000_00010_01000_10000_00000_100110;
RAM[162]<=32'b000000_01101_10000_10000_00000_100110;
RAM[163]<=32'b000000_00101_10000_10000_00000_100110;
//xor reg2 reg3 reg9  reg14 =>reg17
RAM[164]<=32'b000000_00010_00011_10001_00000_100110;
RAM[165]<=32'b000000_01001_10001_10001_00000_100110;
RAM[166]<=32'b000000_01110_10001_10001_00000_100110;
//xor reg11 reg3 reg4 reg10 =>reg18
RAM[167]<=32'b000000_01011_00011_10010_00000_100110;
RAM[168]<=32'b000000_00100_10010_10010_00000_100110;
RAM[169]<=32'b000000_01010_10010_10010_00000_100110;
//��ǰ��+1
RAM[170]<=32'b001000_11010_11010_00000_000000001_00; //addi �����ַreg26+1��reg26
//wb
RAM[171]<=32'b101011_11011_01111_00000_000000000_00; //sw data[reg27+0)   reg15
RAM[172]<=32'b101011_11011_10000_00000_000000100_00; //sw data[reg27+4)   reg16
RAM[173]<=32'b101011_11011_10001_00000_000001000_00; //sw data[reg27+8)   reg17
RAM[174]<=32'b101011_11011_10010_00000_000001100_00; //sw data[reg27+12)  reg18
//ѭ����ת
RAM[175]<=32'b001000_11011_11011_00000_000000001_00; //addi �����ַreg27+1��reg27
RAM[176]<=32'b000101_11010_11111_11111_111010001_00; //bne ���reg26������reg31����������?
//Addroundkey(use reg20 reg21 reg22 reg 23 reg24,fuse reg25)
RAM[177]<=32'b100011_00000_10100_00000_111000011_00; //lw data[451).initial=275->reg20
RAM[178]<=32'b100011_00000_10101_00000_100000010_00; //lw data[258)=259->reg21
RAM[179]<=32'b001000_10101_11001_00000_000010000_00; //addi 259+16 =275->reg25
RAM[180]<=32'b001000_10101_11110_00000_000000001_00; //addi copy to 11110
RAM[181]<=32'b100011_10100_10110_00000_000000000_00; //lw 
RAM[182]<=32'b100011_10101_10000_00000_000000000_00; //lw
RAM[183]<=32'b000000_10110_10000_10001_00000_100110; //xor
RAM[184]<=32'b101011_10101_10001_00000_000000000_00; //sw
RAM[185]<=32'b001000_10100_10100_00000_000000001_00; //addi
RAM[186]<=32'b001000_10101_10101_00000_000000001_00; //addi
RAM[187]<=32'b000101_11110_11001_11111_111111000_00; //bne reg21==reg25? continue:pc-7*4
RAM[188]<=32'b101011_00000_10100_00000_111000011_00; //sw reg20->data[451)
//the BIGround bne end
RAM[189]<=32'b000101_11000_10111_11111_110011100_00; //bne reg23==reg24? continue:pc-99*4











 end
  
 
  
endmodule




module Data_memory(clk,reset,   addr,  we,re ,wdata,rdata);
    //we:write
    //re:read 1=function
    //addr: the high 30 bit is the addr for word (4 byte)
    input   clk, we,re;
    input reset;
    input[31:0]   addr, wdata;
    output[31:0]  rdata; 
    reg[31:0]   RAM[512:0]; 

    //if read, get the data. 
    assign rdata = re ? RAM[addr[31:2]]:0;
    
    //if reset=0 do the reset
    always@(posedge clk or negedge reset)
	 begin
		if (~reset)
		begin
RAM[0]<=32'h63;
RAM[1]<=32'h7c;
RAM[2]<=32'h77;
RAM[3]<=32'h7b;
RAM[4]<=32'hf2;
RAM[5]<=32'h6b;
RAM[6]<=32'h6f;
RAM[7]<=32'hc5;
RAM[8]<=32'h30;
RAM[9]<=32'h01;
RAM[10]<=32'h67;
RAM[11]<=32'h2b;
RAM[12]<=32'hfe;
RAM[13]<=32'hd7;
RAM[14]<=32'hab;
RAM[15]<=32'h76;
RAM[16]<=32'hca;
RAM[17]<=32'h82;
RAM[18]<=32'hc9;
RAM[19]<=32'h7d;
RAM[20]<=32'hfa;
RAM[21]<=32'h59;
RAM[22]<=32'h47;
RAM[23]<=32'hf0;
RAM[24]<=32'had;
RAM[25]<=32'hd4;
RAM[26]<=32'ha2;
RAM[27]<=32'haf;
RAM[28]<=32'h9c;
RAM[29]<=32'ha4;
RAM[30]<=32'h72;
RAM[31]<=32'hc0;
RAM[32]<=32'hb7;
RAM[33]<=32'hfd;
RAM[34]<=32'h93;
RAM[35]<=32'h26;
RAM[36]<=32'h36;
RAM[37]<=32'h3f;
RAM[38]<=32'hf7;
RAM[39]<=32'hcc;
RAM[40]<=32'h34;
RAM[41]<=32'ha5;
RAM[42]<=32'he5;
RAM[43]<=32'hf1;
RAM[44]<=32'h71;
RAM[45]<=32'hd8;
RAM[46]<=32'h31;
RAM[47]<=32'h15;
RAM[48]<=32'h04;
RAM[49]<=32'hc7;
RAM[50]<=32'h23;
RAM[51]<=32'hc3;
RAM[52]<=32'h18;
RAM[53]<=32'h96;
RAM[54]<=32'h05;
RAM[55]<=32'h9a;
RAM[56]<=32'h07;
RAM[57]<=32'h12;
RAM[58]<=32'h80;
RAM[59]<=32'he2;
RAM[60]<=32'heb;
RAM[61]<=32'h27;
RAM[62]<=32'hb2;
RAM[63]<=32'h75;
RAM[64]<=32'h09;
RAM[65]<=32'h83;
RAM[66]<=32'h2c;
RAM[67]<=32'h1a;
RAM[68]<=32'h1b;
RAM[69]<=32'h6e;
RAM[70]<=32'h5a;
RAM[71]<=32'ha0;
RAM[72]<=32'h52;
RAM[73]<=32'h3b;
RAM[74]<=32'hd6;
RAM[75]<=32'hb3;
RAM[76]<=32'h29;
RAM[77]<=32'he3;
RAM[78]<=32'h2f;
RAM[79]<=32'h84;
RAM[80]<=32'h53;
RAM[81]<=32'hd1;
RAM[82]<=32'h00;
RAM[83]<=32'hed;
RAM[84]<=32'h20;
RAM[85]<=32'hfc;
RAM[86]<=32'hb1;
RAM[87]<=32'h5b;
RAM[88]<=32'h6a;
RAM[89]<=32'hcb;
RAM[90]<=32'hbe;
RAM[91]<=32'h39;
RAM[92]<=32'h4a;
RAM[93]<=32'h4c;
RAM[94]<=32'h58;
RAM[95]<=32'hcf;
RAM[96]<=32'hd0;
RAM[97]<=32'hef;
RAM[98]<=32'haa;
RAM[99]<=32'hfb;
RAM[100]<=32'h43;
RAM[101]<=32'h4d;
RAM[102]<=32'h33;
RAM[103]<=32'h85;
RAM[104]<=32'h45;
RAM[105]<=32'hf9;
RAM[106]<=32'h02;
RAM[107]<=32'h7f;
RAM[108]<=32'h50;
RAM[109]<=32'h3c;
RAM[110]<=32'h9f;
RAM[111]<=32'ha8;
RAM[112]<=32'h51;
RAM[113]<=32'ha3;
RAM[114]<=32'h40;
RAM[115]<=32'h8f;
RAM[116]<=32'h92;
RAM[117]<=32'h9d;
RAM[118]<=32'h38;
RAM[119]<=32'hf5;
RAM[120]<=32'hbc;
RAM[121]<=32'hb6;
RAM[122]<=32'hda;
RAM[123]<=32'h21;
RAM[124]<=32'h10;
RAM[125]<=32'hff;
RAM[126]<=32'hf3;
RAM[127]<=32'hd2;
RAM[128]<=32'hcd;
RAM[129]<=32'h0c;
RAM[130]<=32'h13;
RAM[131]<=32'hec;
RAM[132]<=32'h5f;
RAM[133]<=32'h97;
RAM[134]<=32'h44;
RAM[135]<=32'h17;
RAM[136]<=32'hc4;
RAM[137]<=32'ha7;
RAM[138]<=32'h7e;
RAM[139]<=32'h3d;
RAM[140]<=32'h64;
RAM[141]<=32'h5d;
RAM[142]<=32'h19;
RAM[143]<=32'h73;
RAM[144]<=32'h60;
RAM[145]<=32'h81;
RAM[146]<=32'h4f;
RAM[147]<=32'hdc;
RAM[148]<=32'h22;
RAM[149]<=32'h2a;
RAM[150]<=32'h90;
RAM[151]<=32'h88;
RAM[152]<=32'h46;
RAM[153]<=32'hee;
RAM[154]<=32'hb8;
RAM[155]<=32'h14;
RAM[156]<=32'hde;
RAM[157]<=32'h5e;
RAM[158]<=32'h0b;
RAM[159]<=32'hdb;
RAM[160]<=32'he0;
RAM[161]<=32'h32;
RAM[162]<=32'h3a;
RAM[163]<=32'h0a;
RAM[164]<=32'h49;
RAM[165]<=32'h06;
RAM[166]<=32'h24;
RAM[167]<=32'h5c;
RAM[168]<=32'hc2;
RAM[169]<=32'hd3;
RAM[170]<=32'hac;
RAM[171]<=32'h62;
RAM[172]<=32'h91;
RAM[173]<=32'h95;
RAM[174]<=32'he4;
RAM[175]<=32'h79;
RAM[176]<=32'he7;
RAM[177]<=32'hc8;
RAM[178]<=32'h37;
RAM[179]<=32'h6d;
RAM[180]<=32'h8d;
RAM[181]<=32'hd5;
RAM[182]<=32'h4e;
RAM[183]<=32'ha9;
RAM[184]<=32'h6c;
RAM[185]<=32'h56;
RAM[186]<=32'hf4;
RAM[187]<=32'hea;
RAM[188]<=32'h65;
RAM[189]<=32'h7a;
RAM[190]<=32'hae;
RAM[191]<=32'h08;
RAM[192]<=32'hba;
RAM[193]<=32'h78;
RAM[194]<=32'h25;
RAM[195]<=32'h2e;
RAM[196]<=32'h1c;
RAM[197]<=32'ha6;
RAM[198]<=32'hb4;
RAM[199]<=32'hc6;
RAM[200]<=32'he8;
RAM[201]<=32'hdd;
RAM[202]<=32'h74;
RAM[203]<=32'h1f;
RAM[204]<=32'h4b;
RAM[205]<=32'hbd;
RAM[206]<=32'h8b;
RAM[207]<=32'h8a;
RAM[208]<=32'h70;
RAM[209]<=32'h3e;
RAM[210]<=32'hb5;
RAM[211]<=32'h66;
RAM[212]<=32'h48;
RAM[213]<=32'h03;
RAM[214]<=32'hf6;
RAM[215]<=32'h0e;
RAM[216]<=32'h61;
RAM[217]<=32'h35;
RAM[218]<=32'h57;
RAM[219]<=32'hb9;
RAM[220]<=32'h86;
RAM[221]<=32'hc1;
RAM[222]<=32'h1d;
RAM[223]<=32'h9e;
RAM[224]<=32'he1;
RAM[225]<=32'hf8;
RAM[226]<=32'h98;
RAM[227]<=32'h11;
RAM[228]<=32'h69;
RAM[229]<=32'hd9;
RAM[230]<=32'h8e;
RAM[231]<=32'h94;
RAM[232]<=32'h9b;
RAM[233]<=32'h1e;
RAM[234]<=32'h87;
RAM[235]<=32'he9;
RAM[236]<=32'hce;
RAM[237]<=32'h55;
RAM[238]<=32'h28;
RAM[239]<=32'hdf;
RAM[240]<=32'h8c;
RAM[241]<=32'ha1;
RAM[242]<=32'h89;
RAM[243]<=32'h0d;
RAM[244]<=32'hbf;
RAM[245]<=32'he6;
RAM[246]<=32'h42;
RAM[247]<=32'h68;
RAM[248]<=32'h41;
RAM[249]<=32'h99;
RAM[250]<=32'h2d;
RAM[251]<=32'h0f;
RAM[252]<=32'hb0;
RAM[253]<=32'h54;
RAM[254]<=32'hbb;
RAM[255]<=32'h16;
RAM[258]<=32'd1036; //data_addr
RAM[259]<=32'h32;
RAM[260]<=32'h88;
RAM[261]<=32'h31;
RAM[262]<=32'he0;
RAM[263]<=32'h43;
RAM[264]<=32'h5a;
RAM[265]<=32'h31;
RAM[266]<=32'h37;
RAM[267]<=32'hf6;
RAM[268]<=32'h30;
RAM[269]<=32'h98;
RAM[270]<=32'h07;
RAM[271]<=32'ha8;
RAM[272]<=32'h8d;
RAM[273]<=32'ha2;
RAM[274]<=32'h34;
//???1
RAM[275]<=32'h2b;
RAM[276]<=32'h28;
RAM[277]<=32'hab;
RAM[278]<=32'h09;
RAM[279]<=32'h7e;
RAM[280]<=32'hae;
RAM[281]<=32'hf7;
RAM[282]<=32'hcf;
RAM[283]<=32'h15;
RAM[284]<=32'hd2;
RAM[285]<=32'h15;
RAM[286]<=32'h4f;
RAM[287]<=32'h16;
RAM[288]<=32'ha6;
RAM[289]<=32'h88;
RAM[290]<=32'h3c;
//???r
/*
RAM[291]<=32'ha0;
RAM[292]<=32'h88;
RAM[293]<=32'h23;
RAM[294]<=32'h2a;
RAM[295]<=32'hfa;
RAM[296]<=32'h54;
RAM[297]<=32'ha3;
RAM[298]<=32'h6c;
RAM[299]<=32'hfe;
RAM[300]<=32'h2c;
RAM[301]<=32'h39;
RAM[302]<=32'h76;
RAM[303]<=32'h17;
RAM[304]<=32'hb1;
RAM[305]<=32'h39;
RAM[306]<=32'h05;
RAM[307]<=32'hf2;
RAM[308]<=32'h7a;
RAM[309]<=32'h59;
RAM[310]<=32'h73;
RAM[311]<=32'hc2;
RAM[312]<=32'h96;
RAM[313]<=32'h35;
RAM[314]<=32'h59;
RAM[315]<=32'h95;
RAM[316]<=32'hb9;
RAM[317]<=32'h80;
RAM[318]<=32'hf6;
RAM[319]<=32'hf2;
RAM[320]<=32'h43;
RAM[321]<=32'h7a;
RAM[322]<=32'h7f;
RAM[323]<=32'h3d;
RAM[324]<=32'h47;
RAM[325]<=32'h1e;
RAM[326]<=32'h6d;
RAM[327]<=32'h80;
RAM[328]<=32'h16;
RAM[329]<=32'h23;
RAM[330]<=32'h7a;
RAM[331]<=32'h47;
RAM[332]<=32'hfe;
RAM[333]<=32'h7e;
RAM[334]<=32'h88;
RAM[335]<=32'h7d;
RAM[336]<=32'h3e;
RAM[337]<=32'h44;
RAM[338]<=32'h3b;
RAM[339]<=32'hef;
RAM[340]<=32'ha8;
RAM[341]<=32'hb6;
RAM[342]<=32'hdb;
RAM[343]<=32'h44;
RAM[344]<=32'h52;
RAM[345]<=32'h71;
RAM[346]<=32'h0b;
RAM[347]<=32'ha5;
RAM[348]<=32'h5b;
RAM[349]<=32'h25;
RAM[350]<=32'had;
RAM[351]<=32'h41;
RAM[352]<=32'h7f;
RAM[353]<=32'h3b;
RAM[354]<=32'h00;
RAM[355]<=32'hd4;
RAM[356]<=32'h7c;
RAM[357]<=32'hca;
RAM[358]<=32'h11;
RAM[359]<=32'hd1;
RAM[360]<=32'h83;
RAM[361]<=32'hf2;
RAM[362]<=32'hf9;
RAM[363]<=32'hc6;
RAM[364]<=32'h9d;
RAM[365]<=32'hb8;
RAM[366]<=32'h15;
RAM[367]<=32'hf8;
RAM[368]<=32'h87;
RAM[369]<=32'hbc;
RAM[370]<=32'hbc;
RAM[371]<=32'h6d;
RAM[372]<=32'h11;
RAM[373]<=32'hdb;
RAM[374]<=32'hca;
RAM[375]<=32'h88;
RAM[376]<=32'h0b;
RAM[377]<=32'hf9;
RAM[378]<=32'h00;
RAM[379]<=32'ha3;
RAM[380]<=32'h3e;
RAM[381]<=32'h86;
RAM[382]<=32'h93;
RAM[383]<=32'h7a;
RAM[384]<=32'hfd;
RAM[385]<=32'h41;
RAM[386]<=32'hfd;
RAM[387]<=32'h4e;
RAM[388]<=32'h5f;
RAM[389]<=32'h84;
RAM[390]<=32'h4e;
RAM[391]<=32'h54;
RAM[392]<=32'h5f;
RAM[393]<=32'ha6;
RAM[394]<=32'ha6;
RAM[395]<=32'hf7;
RAM[396]<=32'hc9;
RAM[397]<=32'h4f;
RAM[398]<=32'hdc;
RAM[399]<=32'h0e;
RAM[400]<=32'hf3;
RAM[401]<=32'hb2;
RAM[402]<=32'h4f;
RAM[403]<=32'hea;
RAM[404]<=32'hb5;
RAM[405]<=32'h31;
RAM[406]<=32'h7f;
RAM[407]<=32'hd2;
RAM[408]<=32'h8d;
RAM[409]<=32'h2b;
RAM[410]<=32'h8d;
RAM[411]<=32'h73;
RAM[412]<=32'hba;
RAM[413]<=32'hf5;
RAM[414]<=32'h29;
RAM[415]<=32'h21;
RAM[416]<=32'hd2;
RAM[417]<=32'h60;
RAM[418]<=32'h2f;
RAM[419]<=32'hac;
RAM[420]<=32'h19;
RAM[421]<=32'h28;
RAM[422]<=32'h57;
RAM[423]<=32'h77;
RAM[424]<=32'hfa;
RAM[425]<=32'hd1;
RAM[426]<=32'h5c;
RAM[427]<=32'h66;
RAM[428]<=32'hdc;
RAM[429]<=32'h29;
RAM[430]<=32'h00;
RAM[431]<=32'hf3;
RAM[432]<=32'h21;
RAM[433]<=32'h41;
RAM[434]<=32'h6e;
RAM[435]<=32'hd0;
RAM[436]<=32'hc9;
RAM[437]<=32'he1;
RAM[438]<=32'hb6;
RAM[439]<=32'h14;
RAM[440]<=32'hee;
RAM[441]<=32'h3f;
RAM[442]<=32'h63;
RAM[443]<=32'hf9;
RAM[444]<=32'h25;
RAM[445]<=32'h0c;
RAM[446]<=32'h0c;
RAM[447]<=32'ha8;
RAM[448]<=32'h89;
RAM[449]<=32'hc8;
RAM[450]<=32'ha6;  */
RAM[451]<=32'd1100;  //???addr 275*4

//rns
RAM[452]<=32'h01; 
RAM[453]<=32'h02; 
RAM[454]<=32'h04; 
RAM[455]<=32'h08; 
RAM[456]<=32'h10; 
RAM[457]<=32'h20; 
RAM[458]<=32'h40; 
RAM[459]<=32'h80; 
RAM[460]<=32'h1b; 
RAM[461]<=32'h36; 
		end
		else begin
			if(we)  
				RAM[addr[31:2]]<= wdata; 
			else
			    RAM[addr[31:2]]<= RAM[addr[31:2]]; 
		end
	 end

    reg[31:0]   watchdog[15:0];
    always @*
    begin
            watchdog[0]=RAM[259];
            watchdog[1]=RAM[260];
            watchdog[2]=RAM[261];
            watchdog[3]=RAM[262];
            
            watchdog[4]=RAM[263];
            watchdog[5]=RAM[264];
            watchdog[6]=RAM[265];
            watchdog[7]=RAM[266];
            
            watchdog[8]=RAM[267];
            watchdog[9]=RAM[268];
            watchdog[10]=RAM[269];
            watchdog[11]=RAM[270];
            
            watchdog[12]=RAM[271];
            watchdog[13]=RAM[272];
            watchdog[14]=RAM[273];
            watchdog[15]=RAM[274];
                        
    
    end	
endmodule
